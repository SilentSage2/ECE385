module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1 
timeprecision 1ns;

// These signals are internal because the processor will be 
// instantiated as a submodule in testbench.
logic Clk = 0;
logic Reset, Run, Continue;
//logic [11:0] LED
logic CE, UB, LB, OE, WE;
logic [19:0] ADDR;
logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7;
logic [15:0] MAR, MDR, PC, IR, S, R0, R1, R2, R3, R4, R5, R6, R7;
logic [11:0] LED;
logic [4:0] State;
wire [15:0] Data;
	
// A counter to count the instances where simulation results
// do no match with expected results
//integer ErrorCnt = 0;
		
// Instantiating the DUT
// Make sure the module and signal names match with those in your design
lab6_toplevel mt(.*);

assign MAR = mt.my_slc.MAR;
assign MDR = mt.my_slc.MDR;
assign IR = mt.my_slc.IR;
assign PC = mt.my_slc.PC;	
assign R0 = mt.my_slc.reg_file_unit.R0_out;
assign R1 = mt.my_slc.reg_file_unit.R1_out;
assign R2 = mt.my_slc.reg_file_unit.R2_out;
assign R3 = mt.my_slc.reg_file_unit.R3_out;
assign R4 = mt.my_slc.reg_file_unit.R4_out;
assign R5 = mt.my_slc.reg_file_unit.R5_out;
assign R6 = mt.my_slc.reg_file_unit.R6_out;
assign R7 = mt.my_slc.reg_file_unit.R7_out;
assign State = mt.my_slc.state_controller.State;

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

// Testing begins here
// The initial block is not synthesizable
// Everything happens sequentially inside an initial block
// as in a software program
initial begin: TEST_VECTORS
Reset = 0;		// Toggle loadB clearA
Continue = 1;
Run = 1;
//S = 8'h1;	// Specify S --load into B
#10 
Reset = 1;
S = 16'h0014;
#10 Run = 0;

#10 Run = 1;
//
#50
S = 16'h0004;
#10 Continue = 0;
#10 Continue = 1;
//
#50
S = 16'h0003;
#10 Continue = 0;
#10 Continue = 1;

#150 Continue = 0; //BR
#10 Continue = 1;

#150 Continue = 0;
#10 Continue = 1;

end

endmodule
