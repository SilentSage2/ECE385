module shift_reg(

                 );
endmodule
