module audio{
             logic input CLK,      
             logic input Reset,    
        
//         audio_interface signals
             logic output AUD_MCLK
				 logic input AUD_BCLK      
				 logic input AUD_ADCDAT    
				 logic output AUD_DACDAT   
				 logic input AUD_DACLRCK   
				 logic input AUD_ADCLRCK   
				 logic output I2C_SDAT     
				 logic output I2C_SCLK     
             };
				 
				 
audio_interface
				 
endmodule
