module cursor(input logic [5:0] X, Y,
						output logic [4:0] cursor_color
					);
	parameter[0:33][19:0] cursor = {
	20'b10000000000000000000,
	20'b11000000000000000000,
	20'b11100000000000000000,
	20'b11110000000000000000,
	20'b11111100000000000000,
	20'b11111110000000000000,
	20'b11111111000000000000,
	20'b11111111100000000000,
	20'b11111111110000000000,
	20'b11111111111000000000,
	20'b11111111111100000000,
	20'b11111111111110000000,
	20'b11111111111111100000,
	20'b11111111111111110000,
	20'b11111111111111111000,
	20'b11111111111111111100,
	20'b11111111111111111110,
	20'b11111111111111111100,
	20'b11111111111111100000,
	20'b11111111111110000000,
	20'b11111111111110000000,
	20'b11111111111110000000,
	20'b11111100111110000000,
	20'b11110000011111000000,
	20'b11000000011111000000,
	20'b00000000001111100000,
	20'b00000000001111100000,
	20'b00000000001111110000,
	20'b00000000000111110000,
	20'b00000000000111110000,
	20'b00000000000011111000,
	20'b00000000000011111000,
	20'b00000000000001100000,
	20'b00000000000000000000
	};
	
assign cursor_color = cursor[Y][6'd19-X] ? 5'h3 : 5'h0; //output color 0 or color black

endmodule

module shoe(input [5:0] X, Y,
				output [4:0] shoe_color);
	parameter [0:1600-1][4:0] shoe = {
	5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h4,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hb,5'hb,5'hc,5'h3,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hb,5'hc,5'hc,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hb,5'hc,5'hc,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hc,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'h3,5'h3,5'h3,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hc,5'h3,5'h3,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'h2,5'h2,5'hb,5'hb,5'hb,5'hc,5'h3,5'h3,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hb,5'hb,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hb,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hc,5'h3,5'h3,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hb,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hb,5'hc,5'hc,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'h3,5'hc,5'hc,5'hc,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'h3,5'hc,5'h3,5'hc,5'h2,5'h2,5'hb,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'h3,5'h3,5'h3,5'h3,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'h3,5'h3,5'h3,5'h3,5'h2,5'h2,5'h2,5'hb,5'hb,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'h2,5'h2,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'h2,5'h2,5'h2,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hc,5'h2,5'h2,5'h2,5'h2,5'hb,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hb,5'h2,5'h2,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'h2,5'h2,5'h2,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hc,5'h2,5'h2,5'h2,5'h2,5'hb,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hb,5'h2,5'h2,5'h2,5'h2,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'h2,5'h2,5'h2,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hc,5'h2,5'h2,5'h2,5'h2,5'hb,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hb,5'h2,5'h2,5'hb,5'hb,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'h2,5'h2,5'h2,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hc,5'h2,5'h2,5'h2,5'h2,5'hb,5'h3,5'h3,5'h2,5'h2,5'h2,5'h2,5'h2,5'hc,5'h3,5'hb,5'h2,5'h2,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'h2,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'h2,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'h3,5'h3,5'h3,5'h3,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'h3,5'h3,5'h3,5'h3,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'hc,5'hc,5'hc,5'hc,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'hc,5'hc,5'hc,5'hc,5'hc,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h2,5'h2,5'h2,5'h2,5'h2,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,
5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4
	
};

assign shoe_color = shoe[Y*40+X];

endmodule




module bomb_sprite(input logic [5:0] X, Y,
						output logic [4:0] bomb_color
					);
	parameter[0:1600-1][4:0] bomb = {

5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h0,5'h0,5'h3,5'h3,5'h1,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h0,5'h0,5'h3,5'h3,5'h1,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h3,5'h3,5'h1,5'h1,5'h0,5'h0,5'h0,5'h0,5'h1,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h3,5'h3,5'h3,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h3,5'h3,5'h3,5'h1,5'h1,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h3,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h0,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h3,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h0,5'h1,5'h1,5'h0,5'h0,5'h2,5'h2,5'h2,5'h3,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h1,5'h1,5'h0,5'h2,5'h2,5'h3,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h0,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h0,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h0,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h1,5'h1,5'h1,5'h1,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h1,5'h1,5'h1,5'h1,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};
assign bomb_color = bomb[Y*40+X];

endmodule


module bombcenter(input logic [5:0] bcenter_X, bcenter_Y,
						output logic [4:0] bombcenter_color
					);
	parameter[0:1600-1][4:0] bcenter = {

5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h6,5'h3,5'h3,5'h3,5'h3,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h3,5'h3,5'h3,5'h3,
5'h4,5'h4,5'h4,5'h4,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,
5'h3,5'h3,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h3,5'h5,5'h4,5'h4,
5'h3,5'h3,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h3,5'h3,5'h6,5'h4,5'h4

};
assign bombcenter_color = bcenter[bcenter_Y*40+bcenter_X];

endmodule


module bleft(input logic [5:0] X, Y,
						output logic [4:0] bleft_color
					);
	parameter[0:1600-1][4:0] bleft = {
5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h0,5'h0,5'h6,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h4,5'h4,5'h5,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h6,5'h5,5'h4,5'h5,5'h6,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h4,5'h4,5'h5,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,
5'h4,5'h4,5'h5,5'h0,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h0,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h0,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h5,5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,
5'h4,5'h5,5'h6,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,
5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h6,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h5,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4

};
assign bleft_color = bleft[Y*40+X];

endmodule


module bright(input logic [5:0] X, Y,
						output logic [4:0] bright_color
					);
	parameter[0:1600-1][4:0] bright = {
5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h0,5'h0,5'h6,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h5,5'h0,5'h0,5'h6,5'h4,5'h5,5'h0,5'h0,5'h6,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h6,5'h5,5'h4,5'h5,5'h6,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h0,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h5,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,
5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h5,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4
	};
assign bright_color = bright[Y*40+X];

endmodule



module bup(input logic [5:0] X, Y,
						output logic [4:0] bup_color
					);
	parameter[0:1600-1][4:0] bup = {
	
5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h5,5'h0,5'h0,5'h6,5'h4,5'h5,5'h0,5'h0,5'h6,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h0,5'h0,5'h5,5'h4,5'h4,5'h6,5'h0,5'h5,5'h4,5'h4,
5'h4,5'h4,5'h5,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h0,5'h0,
5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h4,5'h4,5'h5,5'h0,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,
5'h6,5'h6,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h0,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0
	
	};
assign bup_color = bup[Y*40+X];

endmodule



module blow(input logic [5:0] X, Y,
						output logic [4:0] blow_color
					);
	parameter[0:1600-1][4:0] blow = {
5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h0,5'h0,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h6,5'h6,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,
5'h4,5'h4,5'h5,5'h0,5'h0,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,
5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h6,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,
5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,
5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h0,5'h0,
5'h4,5'h4,5'h6,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h4,5'h5,5'h6,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h5,5'h5,5'h4,5'h4,5'h4,5'h4,5'h6,5'h0,5'h0,5'h0,5'h0,
5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,
5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h6,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,
5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h6,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h6,5'h6,5'h5,5'h5,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,5'h5,5'h5,5'h6,5'h6,5'h5,5'h4,5'h4,5'h4,5'h5,5'h5,
5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h6,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h0,5'h0,5'h6,5'h5,5'h4,5'h4,5'h4,5'h4,
5'h4,5'h4,5'h4,5'h4,5'h5,5'h6,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h5,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h6,5'h4,5'h4,5'h5,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h5,5'h4,5'h4,5'h4,5'h4

	};
assign blow_color = blow[Y*40+X];

endmodule


module brick(input logic [5:0] brick_X, brick_Y,
						output logic [4:0] brick_color
					);
	parameter[0:1600-1][4:0] brick = {
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h2,5'h2,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h2,5'h1,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h1,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,5'h3,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,
5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2
};

assign brick_color = brick[brick_Y*40+brick_X];

endmodule


module wall(input logic [5:0] wall_X, wall_Y,
						output logic [4:0] wall_color
					);
	parameter[0:1600-1][4:0] wall = {

5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h1,5'h1,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h1,5'h1,5'h2,5'h2,
5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h3,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h1,5'h1,5'h2,5'h2,
5'h1,5'h1,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h1,5'h2,5'h2,5'h2,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,
5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2
};

assign wall_color = wall[wall_Y*40+wall_X];

endmodule

// player1 sprites (front left right back)

module player1_front(input logic [5:0] player1_X, player1_Y,
						output logic [4:0] player1_color
					);
	parameter[0:1600-1][4:0] player1_front = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h11,5'h13,5'h13,5'h11,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h12,5'h12,5'h11,5'h12,5'h11,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h2,5'h12,5'h12,5'h2,5'h11,5'h2,5'h12,5'h11,5'h2,5'h2,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h13,5'h13,5'h12,5'h2,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h2,5'h2,5'h2,5'h2,5'h12,5'h13,5'ha,5'h11,5'h11,5'h2,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h12,5'h11,5'h11,5'h11,5'h3,5'ha,5'h11,5'h11,5'h12,5'h12,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h13,5'h12,5'h13,5'h13,5'h11,5'h13,5'h3,5'h3,5'h11,5'h11,5'h13,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h12,5'h13,5'ha,5'ha,5'h3,5'h3,5'h3,5'ha,5'h13,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h11,5'h2,5'h12,5'h12,5'h13,5'h13,5'h13,5'h13,5'h13,5'h11,5'h12,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h13,5'h12,5'h12,5'h12,5'h12,5'h11,5'h11,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h11,5'h11,5'h11,5'h3,5'h13,5'h3,5'h13,5'h11,5'h11,5'h11,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h13,5'h11,5'h3,5'h3,5'h13,5'h3,5'h3,5'h11,5'h11,5'ha,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h12,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h13,5'h11,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h3,5'h3,5'h11,5'h11,5'h11,5'h13,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h11,5'h3,5'h3,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h13,5'h11,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h13,5'h12,5'h11,5'h11,5'h13,5'h11,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h13,5'h13,5'h11,5'h11,5'h11,5'h12,5'h12,5'h11,5'h11,5'h12,5'h12,5'h11,5'h11,5'h11,5'h13,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h11,5'h12,5'h11,5'h11,5'h11,5'h3,5'h11,5'h11,5'h11,5'h13,5'h11,5'h11,5'h11,5'h12,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h11,5'h11,5'h13,5'h3,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h11,5'h11,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h11,5'h11,5'h13,5'h13,5'h13,5'h13,5'h3,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h3,5'h13,5'h11,5'h11,5'h11,5'h13,5'h3,5'h3,5'h13,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h11,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h11,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h11,5'h11,5'h11,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h13,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h11,5'h13,5'h3,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h13,5'h3,5'h13,5'h13,5'h3,5'h3,5'h3,5'h3,5'h13,5'h3,5'h3,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h3,5'h3,5'h3,5'h3,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player1_color = player1_front[player1_Y*40+player1_X];

endmodule

module player1_left(input logic [5:0] player1_X, player1_Y,
						output logic [4:0] player1_color
					);
	parameter[0:1600-1][4:0] player1_left = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h3,5'h3,5'h11,5'h13,5'h0,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'ha,5'h12,5'h12,5'h12,5'h12,5'h13,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h12,5'h11,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h12,5'h11,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'h2,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h12,5'h2,5'h2,5'h12,5'h11,5'h12,5'h2,5'h12,5'h12,5'h11,5'h12,5'h12,5'h12,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h12,5'h11,5'h12,5'h2,5'h12,5'h12,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h2,5'h12,5'h2,5'h2,5'h13,5'h13,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h2,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h2,5'h2,5'h12,5'h13,5'h13,5'h13,5'h13,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h11,5'ha,5'h11,5'h12,5'h12,5'h13,5'h12,5'h2,5'h12,5'h2,5'h2,5'h12,5'h12,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h13,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h12,5'h2,5'h12,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'ha,5'h3,5'h11,5'h11,5'h13,5'h13,5'h13,5'h12,5'h12,5'h2,5'h12,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h13,5'ha,5'ha,5'ha,5'ha,5'ha,5'h13,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h13,5'h13,5'ha,5'ha,5'h13,5'h11,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h2,5'h2,5'h12,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h13,5'h11,5'h13,5'h11,5'h11,5'h13,5'h11,5'h11,5'h12,5'h2,5'h2,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h11,5'h13,5'h13,5'h11,5'h11,5'h13,5'h13,5'h11,5'h11,5'h12,5'h2,5'h11,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h12,5'h13,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h2,5'h12,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h13,5'h13,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h12,5'h13,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h12,5'h3,5'ha,5'h11,5'h11,5'h11,5'h13,5'h11,5'h11,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h13,5'h13,5'h11,5'h11,5'h11,5'h3,5'ha,5'h11,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h12,5'h11,5'h11,5'h11,5'ha,5'h3,5'h3,5'h11,5'h11,5'h11,5'ha,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'ha,5'h13,5'h11,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h13,5'h11,5'h11,5'h11,5'h13,5'h11,5'h13,5'h11,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h13,5'ha,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h13,5'h11,5'h11,5'h11,5'h12,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h11,5'h11,5'h13,5'h13,5'h13,5'h11,5'h11,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h13,5'ha,5'h11,5'h11,5'ha,5'h3,5'h3,5'h3,5'h3,5'ha,5'h11,5'h11,5'h3,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h13,5'h3,5'h13,5'h13,5'h3,5'h3,5'h3,5'h3,5'ha,5'ha,5'h11,5'h12,5'h13,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h13,5'h3,5'ha,5'ha,5'h3,5'h0,5'h3,5'h3,5'h3,5'h3,5'h11,5'h12,5'ha,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h11,5'ha,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h0,5'h3,5'ha,5'h13,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h13,5'ha,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h13,5'h13,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h13,5'h13,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h13,5'ha,5'h13,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'ha,5'h3,5'h3,5'h3,5'h3,5'h13,5'h13,5'ha,5'ha,5'h13,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h13,5'h3,5'h3,5'h3,5'h3,5'ha,5'h11,5'h11,5'h11,5'h3,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h13,5'h13,5'h13,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player1_color = player1_left[player1_Y*40+player1_X];

endmodule

module player1_right(input logic [5:0] player1_X, player1_Y,
						output logic [4:0] player1_color
					);
	parameter[0:1600-1][4:0] player1_right = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h3,5'h13,5'h11,5'h11,5'h3,5'h13,5'h13,5'h13,5'ha,5'h3,5'h0,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h12,5'h12,5'h12,5'h11,5'h2,5'h2,5'h2,5'h12,5'h11,5'h13,5'h13,5'ha,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h11,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h11,5'ha,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h11,5'h12,5'h12,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h2,5'h12,5'h11,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h12,5'h11,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h2,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h2,5'h12,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'h12,5'h12,5'h11,5'h11,5'h2,5'h2,5'h2,5'h2,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h11,5'h12,5'h11,5'h12,5'h2,5'h12,5'h2,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h2,5'h2,5'h12,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h11,5'h12,5'h11,5'h12,5'h13,5'h13,5'h11,5'h3,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h11,5'h13,5'h13,5'h11,5'h11,5'h3,5'ha,5'ha,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h13,5'ha,5'ha,5'h13,5'h13,5'h3,5'h13,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h13,5'ha,5'ha,5'ha,5'ha,5'h11,5'h13,5'h0,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h11,5'h11,5'h11,5'h13,5'h13,5'h11,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h2,5'h12,5'h2,5'h2,5'h12,5'h11,5'h13,5'h11,5'h11,5'h11,5'h12,5'h13,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'ha,5'h12,5'h2,5'h2,5'h12,5'h11,5'h13,5'h13,5'h11,5'h11,5'ha,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h2,5'h12,5'h11,5'h13,5'h13,5'h13,5'h11,5'h11,5'h11,5'h13,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h11,5'h2,5'h12,5'h11,5'h11,5'h11,5'h13,5'h13,5'h11,5'h13,5'h11,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h12,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h13,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h11,5'h13,5'h13,5'h11,5'h11,5'h11,5'h13,5'ha,5'h11,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h3,5'h3,5'h13,5'h11,5'h11,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h11,5'h11,5'h11,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h13,5'h11,5'h13,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h13,5'h11,5'h11,5'h11,5'ha,5'h11,5'h11,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h11,5'h11,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h11,5'h11,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h11,5'ha,5'h3,5'ha,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'ha,5'ha,5'h3,5'h3,5'h3,5'h3,5'h13,5'h11,5'ha,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h13,5'ha,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h13,5'h3,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h13,5'ha,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h11,5'h11,5'h13,5'ha,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h11,5'h13,5'h13,5'h13,5'ha,5'h3,5'h0,5'h3,5'h3,5'h3,5'h3,5'h13,5'h13,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h11,5'ha,5'h13,5'h13,5'h13,5'ha,5'h3,5'h3,5'h3,5'h3,5'ha,5'h13,5'h11,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h11,5'h13,5'h3,5'ha,5'ha,5'h3,5'h3,5'h3,5'h3,5'h11,5'h11,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h11,5'h12,5'h11,5'h11,5'ha,5'ha,5'h13,5'h11,5'h11,5'h11,5'h13,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h13,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player1_color = player1_right[player1_Y*40+player1_X];

endmodule


module player1_back(input logic [5:0] player1_X, player1_Y,
						output logic [4:0] player1_color
					);
	parameter[0:1600-1][4:0] player1_back = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h13,5'h12,5'h2,5'h12,5'h12,5'h11,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h11,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'h12,5'h12,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h11,5'h12,5'h2,5'h12,5'h12,5'h2,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h11,5'h11,5'h12,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h12,5'h12,5'h11,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h12,5'h12,5'h12,5'h11,5'h12,5'h12,5'h11,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h2,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h2,5'h12,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h2,5'h2,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h12,5'h2,5'h2,5'h2,5'h11,5'h11,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h11,5'h11,5'h11,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h11,5'h11,5'h12,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h11,5'h13,5'h11,5'h11,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h11,5'h11,5'h13,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h13,5'h3,5'h11,5'h11,5'h12,5'h11,5'h13,5'h12,5'h2,5'h12,5'h13,5'h12,5'h12,5'h11,5'h13,5'h3,5'h13,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h3,5'h3,5'h13,5'h11,5'h11,5'h13,5'h13,5'h11,5'h12,5'h11,5'h13,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h3,5'h3,5'h13,5'h12,5'h11,5'h13,5'h13,5'h13,5'h13,5'h11,5'h13,5'h11,5'h11,5'h11,5'h13,5'h3,5'h13,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'ha,5'h11,5'h12,5'h11,5'h13,5'h13,5'h13,5'h11,5'h13,5'h13,5'h13,5'h11,5'h11,5'h13,5'h13,5'h12,5'h11,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h13,5'h13,5'h11,5'h11,5'h13,5'h13,5'h13,5'h11,5'h12,5'h11,5'h11,5'h11,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h11,5'h13,5'h11,5'h11,5'h11,5'h13,5'h11,5'h13,5'h13,5'h13,5'h11,5'h11,5'h11,5'h13,5'h11,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h3,5'h3,5'ha,5'h11,5'h11,5'h11,5'h13,5'h13,5'h13,5'h13,5'h13,5'h11,5'h11,5'h11,5'ha,5'h3,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'ha,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'ha,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'ha,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h11,5'h3,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h13,5'h3,5'ha,5'h13,5'h13,5'h13,5'h13,5'h13,5'h3,5'h3,5'h11,5'h13,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h11,5'ha,5'h3,5'h0,5'h0,5'h3,5'h3,5'h0,5'h0,5'h3,5'ha,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'ha,5'h11,5'h11,5'h3,5'h0,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'ha,5'h13,5'h11,5'h11,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h11,5'h13,5'h3,5'h0,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h11,5'h11,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h11,5'ha,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h3,5'h13,5'h13,5'h13,5'h13,5'h11,5'h11,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h11,5'h12,5'h11,5'ha,5'ha,5'h3,5'h3,5'h3,5'h3,5'h0,5'h3,5'h13,5'ha,5'ha,5'h11,5'h12,5'h13,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h13,5'h11,5'h12,5'h11,5'h13,5'ha,5'h3,5'h3,5'h3,5'ha,5'h13,5'h11,5'h12,5'h11,5'h13,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h11,5'h12,5'h11,5'h11,5'h11,5'h11,5'h11,5'h12,5'h11,5'ha,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h13,5'h13,5'h13,5'h13,5'h13,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player1_color = player1_back[player1_Y*40+player1_X];

endmodule

// player2 sprites (front left right back)

module player2_front(input logic [5:0] player2_X, player2_Y,
						output logic [4:0] player2_color
					);
	parameter[0:1600-1][4:0] player2_front = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h3,5'h14,5'h14,5'h0,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h14,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h14,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h2,5'h2,5'h12,5'h13,5'h14,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h2,5'h2,5'h14,5'ha,5'h13,5'h13,5'h12,5'h14,5'h13,5'h12,5'h14,5'h12,5'h2,5'h2,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h2,5'h14,5'h14,5'h14,5'h13,5'ha,5'ha,5'h13,5'h12,5'h12,5'h12,5'h2,5'h2,5'h14,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'ha,5'h3,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h14,5'h12,5'h12,5'h14,5'h12,5'h12,5'ha,5'h3,5'h12,5'h12,5'h14,5'h12,5'h12,5'h14,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h3,5'h14,5'h14,5'ha,5'h12,5'h13,5'h3,5'h3,5'h13,5'h12,5'h13,5'h13,5'h14,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h13,5'ha,5'ha,5'ha,5'ha,5'ha,5'ha,5'h13,5'h12,5'h12,5'ha,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h3,5'h14,5'h14,5'h14,5'h14,5'h14,5'h13,5'h13,5'h13,5'h13,5'h13,5'h12,5'h12,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'h13,5'h14,5'h14,5'h13,5'h14,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h3,5'h14,5'h3,5'h14,5'h14,5'h3,5'ha,5'ha,5'h3,5'h12,5'h12,5'h12,5'h14,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h3,5'h14,5'h14,5'h14,5'h14,5'h14,5'h3,5'h3,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h14,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h3,5'h14,5'ha,5'h12,5'h14,5'h14,5'h3,5'ha,5'h14,5'h12,5'h14,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'ha,5'h3,5'h12,5'h14,5'h14,5'ha,5'h14,5'h12,5'h14,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h14,5'h3,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h3,5'h14,5'h2,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h2,5'h14,5'h3,5'ha,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h14,5'h12,5'h2,5'h2,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'h14,5'h12,5'h12,5'h2,5'h12,5'h14,5'h14,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h14,5'h12,5'h12,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h14,5'h12,5'h13,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h3,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h3,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'ha,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h14,5'h3,5'ha,5'h14,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h12,5'h14,5'h14,5'h0,5'h0,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h0,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h12,5'h12,5'h14,5'h12,5'h14,5'h12,5'h12,5'h12,5'h14,5'ha,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h3,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h3,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h13,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h13,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'ha,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h14,5'h14,5'h3,5'h3,5'h13,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player2_color = player2_front[player2_Y*40+player2_X];

endmodule

module player2_left(input logic [5:0] player2_X, player2_Y,
						output logic [4:0] player2_color
					);
	parameter[0:1600-1][4:0] player2_left = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h14,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h13,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h13,5'h13,5'h13,5'h13,5'h13,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'ha,5'h14,5'h12,5'h12,5'h14,5'h13,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'ha,5'h14,5'h12,5'h14,5'h12,5'h13,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h14,5'h14,5'h12,5'h14,5'h13,5'ha,5'h14,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'ha,5'ha,5'h13,5'ha,5'ha,5'ha,5'h13,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h14,5'ha,5'ha,5'ha,5'ha,5'h13,5'h12,5'h12,5'h2,5'h14,5'h12,5'h2,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h2,5'h14,5'h12,5'h2,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h13,5'ha,5'h12,5'h12,5'h12,5'h12,5'h2,5'h14,5'h3,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h13,5'h12,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h3,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h12,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h2,5'h14,5'ha,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h2,5'h14,5'ha,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h14,5'h14,5'h14,5'h12,5'h2,5'h12,5'h14,5'h14,5'h14,5'h2,5'h14,5'h0,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'ha,5'h14,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h12,5'ha,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h2,5'h14,5'h14,5'h12,5'h12,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h12,5'h2,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h2,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h13,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'h2,5'h14,5'h14,5'h14,5'h2,5'h2,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h14,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'ha,5'h3,5'h14,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h13,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'h12,5'h14,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player2_color = player2_left[player2_Y*40+player2_X];

endmodule

module player2_right(input logic [5:0] player2_X, player2_Y,
						output logic [4:0] player2_color
					);
	parameter[0:1600-1][4:0] player2_right = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'ha,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'h13,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h13,5'h14,5'h14,5'h13,5'ha,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h14,5'h13,5'h12,5'h12,5'h12,5'ha,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h13,5'h14,5'h14,5'h12,5'h12,5'h14,5'h13,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'ha,5'h13,5'h13,5'h12,5'h12,5'h14,5'ha,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'ha,5'h14,5'h14,5'ha,5'ha,5'ha,5'h13,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h2,5'h14,5'h2,5'h12,5'h12,5'h14,5'h13,5'ha,5'ha,5'h13,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h2,5'h12,5'ha,5'h12,5'h12,5'h14,5'h13,5'h14,5'h14,5'h14,5'h12,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h14,5'h14,5'h12,5'h12,5'h12,5'h13,5'h14,5'h3,5'h3,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h14,5'h3,5'h12,5'ha,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h3,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h13,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h14,5'h0,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h14,5'h13,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h0,5'h12,5'h14,5'h14,5'h14,5'ha,5'h12,5'h14,5'h12,5'h12,5'h14,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h0,5'h3,5'h12,5'h14,5'h14,5'ha,5'h14,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h14,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'ha,5'h14,5'h12,5'h12,5'h12,5'h14,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h14,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h2,5'h14,5'h12,5'h2,5'h2,5'h12,5'h14,5'h14,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h14,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h2,5'h12,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h14,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h14,5'h12,5'h2,5'h12,5'h12,5'h2,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h14,5'ha,5'h14,5'h14,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player2_color = player2_right[player2_Y*40+player2_X];

endmodule


module player2_back(input logic [5:0] player2_X, player2_Y,
						output logic [4:0] player2_color
					);
	parameter[0:1600-1][4:0] player2_back = {


5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h2,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h2,5'h2,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h12,5'h2,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h12,5'h12,5'h2,5'h2,5'h12,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h2,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h2,5'h12,5'ha,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h2,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h2,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h12,5'h12,5'h12,5'h2,5'h2,5'h2,5'h12,5'h12,5'h2,5'h2,5'h2,5'h14,5'h14,5'h14,5'h3,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h14,5'h14,5'h12,5'h2,5'h2,5'h2,5'h2,5'h2,5'h12,5'h14,5'h3,5'h3,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h2,5'h14,5'h14,5'h12,5'h2,5'h12,5'h12,5'h2,5'h2,5'h14,5'h14,5'h3,5'h3,5'h3,5'h3,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h12,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h12,5'h12,5'h3,5'h3,5'h14,5'h14,5'h3,5'h3,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'h12,5'h14,5'h2,5'h12,5'h14,5'h12,5'h12,5'h14,5'h3,5'h3,5'h14,5'h12,5'h3,5'h3,5'h3,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'ha,5'h14,5'h14,5'h12,5'h2,5'h12,5'h14,5'h12,5'h12,5'h12,5'ha,5'h3,5'h3,5'h12,5'h14,5'h3,5'ha,5'ha,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'h14,5'ha,5'h14,5'h2,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h12,5'h12,5'ha,5'h12,5'h12,5'h14,5'h14,5'h3,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h14,5'h14,5'h12,5'h2,5'h2,5'h12,5'h14,5'h12,5'h14,5'h14,5'h14,5'h12,5'h2,5'h2,5'h2,5'h12,5'h14,5'h12,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'ha,5'h12,5'h13,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h12,5'h12,5'h13,5'h12,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h14,5'ha,5'h12,5'h12,5'h14,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h12,5'h14,5'h13,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h3,5'h14,5'ha,5'h0,5'h12,5'h2,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h2,5'h14,5'h0,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h2,5'h12,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h2,5'h14,5'h14,5'h12,5'h14,5'h14,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h14,5'h14,5'h14,5'h12,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h12,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h12,5'h14,5'h12,5'h2,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h14,5'h12,5'h14,5'h14,5'h12,5'h14,5'h12,5'h2,5'h12,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'h14,5'h12,5'h12,5'h12,5'h12,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h14,5'h14,5'h14,5'h13,5'h0,5'h0,5'h14,5'h14,5'h14,5'h14,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};

assign player2_color = player2_back[player2_Y*40+player2_X];

endmodule

// treasure sprites (hat and liquid)

module hat(input logic [5:0] X, Y,
						output logic [4:0] hat_color
					);
	parameter[0:1600-1][4:0] hat = {
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h0,5'h10,5'h10,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'hf,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'hf,5'h0,5'hf,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h10,5'h0,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h10,5'h0,5'h0,5'hf,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'hf,5'hf,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'hf,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'hf,5'hf,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'hf,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'hf,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'hf,5'h10,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'h0,5'h10,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h10,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'hf,5'h10,5'h0,5'h0,5'h10,5'h10,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'hf,5'hf,5'hf,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'hf,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'hf,5'h10,5'h10,5'hf,5'hf,5'h10,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'hf,5'h0,5'h0,5'h0,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h0,5'h0,5'h0,5'h0,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hf,5'h10,5'h10,5'h10,5'h10,5'hf,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h10,5'h10,5'h10,5'h10,5'h10,5'h10,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0

	};
assign hat_color = hat[Y*40+X];

endmodule


module liquid(input logic [5:0] X, Y,
						output logic [4:0] liquid_color
					);
	parameter[0:1600-1][4:0] liquid = {

5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'he,5'he,5'he,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'he,5'he,5'he,5'he,5'he,5'he,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'hd,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'hd,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'hc,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'hd,5'hd,5'hc,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'hb,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'h0,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'he,5'he,5'he,5'he,5'he,5'he,5'he,5'hd,5'h0,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'he,5'he,5'he,5'he,5'he,5'hd,5'h0,5'hd,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hc,5'he,5'he,5'hc,5'h0,5'h0,5'hd,5'hc,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hd,5'hc,5'hd,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hd,5'hd,5'hc,5'hc,5'hd,5'hc,5'hc,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hc,5'hc,5'hd,5'hc,5'hc,5'hc,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hc,5'hc,5'hc,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hd,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hc,5'hd,5'hc,5'hb,5'hc,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hd,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hc,5'hd,5'hc,5'hc,5'hb,5'hc,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'h0,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hd,5'hc,5'hb,5'hc,5'hb,5'hc,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hd,5'hd,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'hc,5'hb,5'hc,5'hc,5'hb,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hb,5'hb,5'hc,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hc,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hb,5'hb,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hb,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hc,5'hc,5'hc,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hb,5'hc,5'hc,5'hc,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hc,5'hd,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'hd,5'hd,5'hd,5'hd,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,
5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0,5'h0
};
assign liquid_color = liquid[Y*40+X];

endmodule




