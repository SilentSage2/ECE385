module multipilication(
                       input [7:0] A,
							  input [7:0] B,
							  output [15:0] Product,
							  output CO
							  );
							  
endmodule	