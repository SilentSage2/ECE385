module startpage(
				input logic Clk,
				input logic load_startpage,
				